//Pipeline Controller skeleton
//TODOS:
//add logic, add outputs needed that were added to Project2.v for the pipeline processor
module PipelineController(EX_op, EX_func, MEM_op, MEM_func, WB_op, WB_func, 
								  allowBr, brBaseMux, rs1Mux, rs2Mux, alu2Mux, 
								  aluOp, cmpOp, wrReg, wrMem, dstRegMux);

								  
endmodule								  